LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE MY_PACKAGE IS

COMPONENT Counter IS
	GENERIC	(Ceil_value: INTEGER);

	PORT	(
		Clk, Inc, Clr:	IN STD_LOGIC;
		Z:			OUT STD_LOGIC;
		Count:	OUT INTEGER RANGE 0 TO Ceil_value
		);
END COMPONENT;

COMPONENT Data_out IS
	GENERIC (
		ROW_SIZE:		INTEGER;
		COL_SIZE:		INTEGER
		);
	
	PORT	(
		Clk:		IN STD_LOGIC;
		We_out:	IN STD_LOGIC;
		Re_out:	IN STD_LOGIC;
		Addr:		IN INTEGER RANGE 0 TO ROW_SIZE * COL_SIZE - 1;
		Din:		IN INTEGER;
		Dout:		OUT INTEGER
		);		
END COMPONENT;

COMPONENT Data_in IS
	GENERIC (
		ROW_SIZE:		INTEGER;
		COL_SIZE:		INTEGER
		);
	
	PORT	(
		Clk:		IN STD_LOGIC;
		We_in:	IN STD_LOGIC;
		Re_in:	IN STD_LOGIC;
		Addr:		IN INTEGER RANGE 0 TO ROW_SIZE * COL_SIZE - 1;
		Din:		IN INTEGER;
		Dout:		OUT INTEGER
		);		
END COMPONENT;

COMPONENT Controller IS

	PORT	(
		Start:	IN STD_LOGIC;
		Clk:		IN STD_LOGIC;
		Reset:	IN STD_LOGIC;
		R_z, Rs_z, C_z, Cs_z, Gt:			IN STD_LOGIC;
		R_clr, Rs_Clr, C_clr, Cs_clr:	OUT STD_LOGIC;
		R_inc, Rs_inc, C_inc, Cs_inc:	OUT STD_LOGIC;
		Re_in, Re_out, We_in, We_out:	OUT STD_LOGIC;
		Done:		OUT STD_LOGIC
		);
END COMPONENT;

COMPONENT Datapath IS
	GENERIC	(
		ROW_IN:		INTEGER;
		COL_IN:		INTEGER;
		ROW_OUT:	INTEGER;
		COL_OUT:	INTEGER;
		ROW_STEP:	INTEGER;
		COL_STEP:	INTEGER
		);

	
	PORT	(
		Clk:	IN STD_LOGIC;
		R_clr, Rs_clr, C_clr, Cs_clr:	IN STD_LOGIC;
		R_inc, Rs_inc, C_inc, Cs_inc:	IN STD_LOGIC;
		Data_in, Data_out:	IN INTEGER;
		R_z, Rs_z, C_z, Cs_z, Gt:		OUT STD_LOGIC;
		Data_in_addr:		OUT INTEGER RANGE 0 TO ROW_IN * COL_IN - 1;
		Data_out_addr:	OUT INTEGER RANGE 0 TO ROW_OUT * COL_OUT - 1
		);
END COMPONENT;

COMPONENT Max_pooling IS
	GENERIC	(
		ROW_IN:		INTEGER;
		COL_IN:		INTEGER;
		ROW_OUT:	INTEGER;
		COL_OUT:	INTEGER;
		ROW_STEP:	INTEGER;
		COL_STEP:	INTEGER
		);
		
	PORT	(
		Clk:		IN STD_LOGIC;
		Start:	IN STD_LOGIC;
		Reset:	IN STD_LOGIC;		
		Done:		OUT STD_LOGIC
		);	
END COMPONENT;	

END PACKAGE MY_PACKAGE;

